module prefix_32(s,cout,x,y,cin);
output[31:0]s;
output cout;
input wire[31:0]x,y;
input cin;


wire[31:0]g,a,p;
wire[36:0]g1,a1;
wire[32:0]c;

g_a ga1(g[0],a[0],p[0],x[0],y[0]);
g_a ga2(g[1],a[1],p[1],x[1],y[1]);
g_a ga3(g[2],a[2],p[2],x[2],y[2]);
g_a ga4(g[3],a[3],p[3],x[3],y[3]);
g_a ga5(g[4],a[4],p[4],x[4],y[4]);
g_a ga6(g[5],a[5],p[5],x[5],y[5]);
g_a ga7(g[6],a[6],p[6],x[6],y[6]);
g_a ga8(g[7],a[7],p[7],x[7],y[7]);
g_a ga9(g[8],a[8],p[8],x[8],y[8]);
g_a ga10(g[9],a[9],p[9],x[9],y[9]);
g_a ga11(g[10],a[10],p[10],x[10],y[10]);
g_a ga12(g[11],a[11],p[11],x[11],y[11]);
g_a ga13(g[12],a[12],p[12],x[12],y[12]);
g_a ga14(g[13],a[13],p[13],x[13],y[13]);
g_a ga15(g[14],a[14],p[14],x[14],y[14]);
g_a ga16(g[15],a[15],p[15],x[15],y[15]);
g_a ga17(g[16],a[16],p[16],x[16],y[16]);
g_a ga18(g[17],a[17],p[17],x[17],y[17]);
g_a ga19(g[18],a[18],p[18],x[18],y[18]);
g_a ga20(g[19],a[19],p[19],x[19],y[19]);
g_a ga21(g[20],a[20],p[20],x[20],y[20]);
g_a ga22(g[21],a[21],p[21],x[21],y[21]);
g_a ga23(g[22],a[22],p[22],x[22],y[22]);
g_a ga24(g[23],a[23],p[23],x[23],y[23]);
g_a ga25(g[24],a[24],p[24],x[24],y[24]);
g_a ga26(g[25],a[25],p[25],x[25],y[25]);
g_a ga27(g[26],a[26],p[26],x[26],y[26]);
g_a ga28(g[27],a[27],p[27],x[27],y[27]);
g_a ga29(g[28],a[28],p[28],x[28],y[28]);
g_a ga30(g[29],a[29],p[29],x[29],y[29]);
g_a ga31(g[30],a[30],p[30],x[30],y[30]);
g_a ga32(g[31],a[31],p[31],x[31],y[31]);

dot d1(c[1],g[0],a[0],cin);
circle c1(g1[0],a1[0],g[2],a[2],g[1],a[1]);
circle c2(g1[1],a1[1],g[4],a[4],g[3],a[3]);
circle c3(g1[2],a1[2],g[6],a[6],g[5],a[5]);
circle c4(g1[3],a1[3],g[8],a[8],g[7],a[7]);
circle c5(g1[4],a1[4],g[10],a[10],g[9],a[9]);
circle c6(g1[5],a1[5],g[12],a[12],g[11],a[11]);
circle c7(g1[6],a1[6],g[14],a[14],g[13],a[13]);
circle c8(g1[7],a1[7],g[16],a[16],g[15],a[15]);
circle c9(g1[8],a1[8],g[18],a[18],g[17],a[17]);
circle c10(g1[9],a1[9],g[20],a[20],g[19],a[19]);
circle c11(g1[10],a1[10],g[22],a[22],g[21],a[21]);
circle c12(g1[11],a1[11],g[24],a[24],g[23],a[23]);
circle c13(g1[12],a1[12],g[26],a[26],g[25],a[25]);
circle c14(g1[13],a1[13],g[28],a[28],g[27],a[27]);
circle c15(g1[14],a1[14],g[30],a[30],g[29],a[29]);


dot d2(c[2],g[1],a[1],c[1]);
dot d3(c[3],g1[0],a1[0],c[1]);
circle c16(g1[15],a1[15],g[5],a[5],g1[1],a1[1]);
circle c17(g1[16],a1[16],g1[2],a1[2],g1[1],a1[1]);
circle c18(g1[17],a1[17],g[9],a[9],g1[3],a1[3]);
circle c19(g1[18],a1[18],g1[4],a1[4],g1[3],a1[3]);
circle c20(g1[19],a1[19],g[17],a[17],g1[7],a1[7]);
circle c21(g1[20],a1[20],g1[8],a1[8],g1[7],a1[7]);


dot d4(c[4],g[3],a[3],c[3]);
dot d5(c[5],g1[1],a1[1],c[3]);
dot d6(c[6],g1[7],a1[7],c[3]);
dot d7(c[7],g1[8],a1[8],c[3]);
circle c22(g1[21],a1[21],g[11],a[11],g1[18],a1[18]);
circle c23(g1[22],a1[22],g1[5],a1[5],g1[18],a1[18]);
circle c24(g1[23],a1[23],g[13],a[13],g1[18],a1[18]);
circle c25(g1[24],a1[24],g1[6],a1[6],g1[18],a1[18]);
circle c26(g1[25],a1[25],g[19],a[19],g1[20],a1[20]);
circle c27(g1[26],a1[26],g1[9],a1[9],g1[20],a1[20]);
circle c28(g1[27],a1[27],g[21],a[21],g1[20],a1[20]);
circle c29(g1[28],a1[28],g1[10],a1[10],g1[20],a1[20]);



dot d8(c[8],g[7],a[7],c[7]);
dot d9(c[9],g1[3],a1[3],c[7]);
dot d10(c[10],g1[17],a1[17],c[7]);
dot d11(c[11],g1[18],a1[18],c[7]);
dot d12(c[12],g1[21],a1[21],c[7]);
dot d13(c[13],g1[22],a1[22],c[7]);
dot d14(c[14],g1[23],a1[23],c[7]);
dot d15(c[15],g1[24],a1[24],c[7]);
circle c30(g1[29],a1[29],g[23],a[23],g1[28],a1[28]);
circle c31(g1[30],a1[30],g1[11],a1[11],g1[20],a1[20]);
circle c32(g1[31],a1[31],g[25],a[25],g1[28],a1[28]);
circle c33(g1[32],a1[32],g1[12],a1[12],g1[28],a1[28]);
circle c34(g1[33],a1[33],g[27],a[27],g1[28],a1[28]);
circle c35(g1[34],a1[34],g1[13],a1[13],g1[28],a1[28]);
circle c36(g1[35],a1[35],g[29],a[29],g1[28],a1[28]);
circle c37(g1[36],a1[36],g1[14],a1[14],g1[28],a1[28]);


dot d16(c[16],g[15],a[15],c[15]);
dot d17(c[17],g1[7],a1[7],c[15]);
dot d18(c[18],g1[19],a1[19],c[15]);
dot d19(c[19],g1[20],a1[20],c[15]);
dot d20(c[20],g1[25],a1[25],c[15]);
dot d21(c[21],g1[26],a1[26],c[15]);
dot d22(c[22],g1[27],a1[27],c[15]);
dot d23(c[23],g1[28],a1[28],c[15]);
dot d24(c[24],g1[29],a1[29],c[15]);
dot d25(c[25],g1[30],a1[30],c[15]);
dot d26(c[26],g1[31],a1[31],c[15]);
dot d27(c[27],g1[32],a1[32],c[15]);
dot d28(c[28],g1[33],a1[33],c[15]);
dot d29(c[29],g1[34],a1[34],c[15]);
dot d30(c[30],g1[35],a1[35],c[15]);
dot d31(c[31],g1[36],a1[36],c[15]);



dot d32(cout,g[31],a[31],c[31]);


assign s[0]=p[0]^cin;
assign s[1]=p[1]^c[1];
assign s[2]=p[2]^c[2];
assign s[3]=p[3]^c[3];
assign s[4]=p[4]^c[4];
assign s[5]=p[5]^c[5];
assign s[6]=p[6]^c[6];
assign s[7]=p[7]^c[7];
assign s[8]=p[8]^c[8];
assign s[9]=p[9]^c[9];
assign s[10]=p[10]^c[10];
assign s[11]=p[11]^c[11];
assign s[12]=p[12]^c[12];
assign s[13]=p[13]^c[13];
assign s[14]=p[14]^c[14];
assign s[15]=p[15]^c[15];
assign s[16]=p[16]^c[16];
assign s[17]=p[17]^c[17];
assign s[18]=p[18]^c[18];
assign s[19]=p[19]^c[19];
assign s[20]=p[20]^c[20];
assign s[21]=p[21]^c[21];
assign s[22]=p[22]^c[22];
assign s[23]=p[23]^c[23];
assign s[24]=p[24]^c[24];
assign s[25]=p[25]^c[25];
assign s[26]=p[26]^c[26];
assign s[27]=p[27]^c[27];
assign s[28]=p[28]^c[28];
assign s[29]=p[29]^c[29];
assign s[30]=p[30]^c[30];
assign s[31]=p[31]^c[31];


endmodule






